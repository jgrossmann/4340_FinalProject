class c_514_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_514_12;
    c_514_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz11x0x0z1110z0xzzxxz10xxxx0xx1zzzzzxzzxxzxxxxxxzxxxxzzxxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
