class c_970_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_970_12;
    c_970_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1101zz110101z11z1x0x1x01xx01z1x1zxzzxxxxxxzzxxxxzxzzxxzzxxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
