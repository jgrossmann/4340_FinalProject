module rr_register_1000_test.sv();

  bit clk = 1;
  bit reset;
  bit change_order_i;
  logic [3:0] priority_order_o;

  


endmodule
