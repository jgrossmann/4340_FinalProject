class c_957_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_957_12;
    c_957_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00x1011z01z0z1100x1zzxxxz0xx0x0xzzxxzxzzzzxxxxxzzxxxxzzxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
