class c_708_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_708_12;
    c_708_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1x0z0x001z1xxx1xx01x1zxx00x110xzzzxxzxxzzzzzzzxzxzzxxzxzxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
