class c_733_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_733_12;
    c_733_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx0x01zx0xz010x1z0x0z0z111x11zxzzzzzxxxzxzxxzzzzxzzxzxxzzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
