class c_679_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_679_12;
    c_679_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1101z0z01x1xx1z0z1zzz1xzxz1x1z1zxxxzzxzzxzxzzxxxzxzzzzzzxxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
