class c_182_16;
    integer y_pos = 2;
    integer x_pos = 3;
    rand bit[15:0] l_arb_address_i = 16'h5c25; // rand_mode = OFF 

    constraint c_this    // (constraint_mode = ON) (../arbiter/arbiter_transaction.sv:51)
    {
       ((l_arb_address_i[3:0]) <= 4'h3);
    }
endclass

program p_182_16;
    c_182_16 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001x1x10zz0zz1x00xz11z1xzxx1x1z0xxxxxxzzzxzxxzxxxxxzxxxzzxzzzzzz";
            obj.set_randstate(randState);
            obj.l_arb_address_i.rand_mode(0);
            obj.randomize();
        end
endprogram
