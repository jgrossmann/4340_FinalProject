`include "tb/router_class.sv"
class network;

	router r1;
	router r2;
	router r3;
	router r4;
	router r5;
	router r6;
	router r7;
	router r8;
	router r9;
	router r10;
	router r11;
	router r12;
	router r13;
	router r14;
	router r15;
	router r16;

	function new();
		r1 = new(0, 0);
		r2 = new(0, 1);
		r3 = new(0, 2);
		r4 = new(0, 3);
		r5 = new(1, 0);
		r6 = new(1, 1);
		r7 = new(1, 2);
		r8 = new(1, 3);
		r9 = new(2, 0);
		r10 = new(2, 1);
		r11 = new(2, 2);
		r12 = new(2, 3);
		r13 = new(3, 0);
		r14 = new(3, 1);
		r15 = new(3, 2);
		r16 = new(3, 3);
	
	endfunction


endclass
