class c_568_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_568_12;
    c_568_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0x0zx1x1011x0zxzxx01z1x010x100xzzxxzxxxxzxzzzxzzzzzxxzzzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
