module sw_corner_router
(
	input [15 : 0] n_data_i,
	input [15 : 0] e_data_i,
	input [15 : 0] l_data_i,
	input n_valid_i,
	input e_valid_i,
	input l_valid_i,
	input n_credit_i,
	input e_credit_i,
	input l_credit_i,
	output [15 : 0] n_data_o,
	output [15 : 0] e_data_o,
	output [15 : 0] l_data_o,
	output n_valid_o,
	output e_valid_o,
	output l_valid_o,
	output n_credit_o,
	output e_credit_o,
	output l_credit_o,
	input clk,
	input reset
);

endmodule
