module arbiter();

endmodule
