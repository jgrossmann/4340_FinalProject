class c_430_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_430_12;
    c_430_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z00000zx0x110z1x0x01xx10z1011z1zxxxzxzzxxxxxxxzzzxxxzzzxxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
