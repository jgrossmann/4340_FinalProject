module noc (ifc.dut ifc);

endmodule