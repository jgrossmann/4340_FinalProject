class c_571_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_571_12;
    c_571_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzx1z1x0z1z1x01x11z01xxzz0z01zxxzxzzxzzxzzzxzxzzxxzxzzzzxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
