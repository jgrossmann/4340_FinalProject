class flit;


endclass
