class c_618_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_618_12;
    c_618_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111xz1xxz0z1z101x1z0x0xzzxxx0z0xxzzxzxxxxzxzzxzzzzzxxxxzxzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
