class c_758_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_758_12;
    c_758_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1000x10x0xzz0100z01xzxz10101z0zzxxxxzzzxzxzzzzxxxzxzxxzzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
