class c_327_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_327_12;
    c_327_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10xzx110x0z0x0z1zxz0111z1x1x0x00xzzzzzzxzzxxzzxxxxzxxzxxxzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
