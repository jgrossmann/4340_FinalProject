class arbiter;





endclass