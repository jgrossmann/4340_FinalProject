class c_727_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_727_12;
    c_727_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0x0x0xz0x1x01zzxzz0x0z010zz001zzzzxxxxxxzzxxzzxzzzxzxxxxzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
