class mux;





endclass