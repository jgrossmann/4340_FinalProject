class credit_counter;

	logic credit_count;




endclass