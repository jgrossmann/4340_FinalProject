class input_buffer;





endclass