class c_1051_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_1051_12;
    c_1051_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z000z1x010x0x1z1z0x000x1xz1z010zxzxxxxxxxxzzzxzxxxxzxzzxxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
