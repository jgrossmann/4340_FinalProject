class checker;

endclass