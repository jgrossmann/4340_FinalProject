class c_814_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_814_12;
    c_814_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0111zz0x10zz001110zx0x01x1xz1z1zzxzxxzzxxzzzzxzzzxzzzzzxzxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
