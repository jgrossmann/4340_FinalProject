class c_757_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_757_12;
    c_757_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001z0zx01x0z0x000z11xx0xx0x1z1z0xxxzzzxxxzxzzxxxzxzzzzzxxzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
