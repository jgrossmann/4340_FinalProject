class environment;

endclass