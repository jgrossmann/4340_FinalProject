class c_911_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_911_12;
    c_911_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111xxxz00z010xz0z0xx0zz0xxz0z1x1xxxzxzxxxxxxzzzxzzxxxxzxxzzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
