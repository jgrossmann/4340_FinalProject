class c_569_12;
    integer y_pos = 2060830875;
    rand bit[7:0] n_arb_address_i; // rand_mode = ON 

    constraint c_this    // (constraint_mode = ON) (arbiter_transaction.sv:27)
    {
       ((n_arb_address_i[3:0]) >= y_pos);
    }
endclass

program p_569_12;
    c_569_12 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz0x1zz1zz1x01100011xz10x00z00zxzzxzzzzzzxxzzxxxzzxxzzzzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
