class transaction;





endclass